// Copyright (C) 2023  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// PROGRAM		"Quartus Prime"
// VERSION		"Version 22.1std.2 Build 922 07/20/2023 SC Lite Edition"
// CREATED		"Tue Oct  3 16:21:13 2023"

module HD3(
	Reset,
	Clock,
	Sb,
	Sc,
	Sd,
	Se,
	Sf,
	Sg,
	Sa,
	count3,
	count2,
	count1,
	count0
);


input wire	Reset;
input wire	Clock;
output wire	Sb;
output wire	Sc;
output wire	Sd;
output wire	Se;
output wire	Sf;
output wire	Sg;
output wire	Sa;
output wire	count3;
output wire	count2;
output wire	count1;
output wire	count0;

reg	SYNTHESIZED_WIRE_81;
reg	SYNTHESIZED_WIRE_82;
wire	SYNTHESIZED_WIRE_83;
wire	SYNTHESIZED_WIRE_1;
wire	SYNTHESIZED_WIRE_84;
wire	SYNTHESIZED_WIRE_85;
reg	SYNTHESIZED_WIRE_86;
wire	SYNTHESIZED_WIRE_87;
wire	SYNTHESIZED_WIRE_88;
wire	SYNTHESIZED_WIRE_89;
reg	SYNTHESIZED_WIRE_90;
wire	SYNTHESIZED_WIRE_91;
wire	SYNTHESIZED_WIRE_15;
wire	SYNTHESIZED_WIRE_16;
wire	SYNTHESIZED_WIRE_17;
wire	SYNTHESIZED_WIRE_18;
wire	SYNTHESIZED_WIRE_92;
wire	SYNTHESIZED_WIRE_52;
wire	SYNTHESIZED_WIRE_53;
wire	SYNTHESIZED_WIRE_54;
wire	SYNTHESIZED_WIRE_55;
wire	SYNTHESIZED_WIRE_56;
wire	SYNTHESIZED_WIRE_57;
wire	SYNTHESIZED_WIRE_58;
wire	SYNTHESIZED_WIRE_59;
wire	SYNTHESIZED_WIRE_60;
wire	SYNTHESIZED_WIRE_61;
wire	SYNTHESIZED_WIRE_62;
wire	SYNTHESIZED_WIRE_63;
wire	SYNTHESIZED_WIRE_64;
wire	SYNTHESIZED_WIRE_65;
wire	SYNTHESIZED_WIRE_66;
wire	SYNTHESIZED_WIRE_67;
wire	SYNTHESIZED_WIRE_68;
wire	SYNTHESIZED_WIRE_77;
wire	SYNTHESIZED_WIRE_78;
wire	SYNTHESIZED_WIRE_79;
wire	SYNTHESIZED_WIRE_80;

assign	count3 = SYNTHESIZED_WIRE_90;
assign	count2 = SYNTHESIZED_WIRE_86;
assign	count1 = SYNTHESIZED_WIRE_82;
assign	count0 = SYNTHESIZED_WIRE_81;
assign	SYNTHESIZED_WIRE_84 = 1;



assign	SYNTHESIZED_WIRE_91 =  ~SYNTHESIZED_WIRE_81;

assign	SYNTHESIZED_WIRE_88 =  ~SYNTHESIZED_WIRE_82;


always@(posedge SYNTHESIZED_WIRE_83 or negedge Reset or negedge SYNTHESIZED_WIRE_84)
begin
if (!Reset)
	begin
	SYNTHESIZED_WIRE_81 <= 0;
	end
else
if (!SYNTHESIZED_WIRE_84)
	begin
	SYNTHESIZED_WIRE_81 <= 1;
	end
else
	begin
	SYNTHESIZED_WIRE_81 <= SYNTHESIZED_WIRE_1;
	end
end


always@(posedge Clock or negedge Reset or negedge SYNTHESIZED_WIRE_84)
begin
if (!Reset)
	begin
	SYNTHESIZED_WIRE_90 <= 0;
	end
else
if (!SYNTHESIZED_WIRE_84)
	begin
	SYNTHESIZED_WIRE_90 <= 1;
	end
else
	begin
	SYNTHESIZED_WIRE_90 <= SYNTHESIZED_WIRE_85;
	end
end

assign	SYNTHESIZED_WIRE_18 = SYNTHESIZED_WIRE_81 | SYNTHESIZED_WIRE_86 | SYNTHESIZED_WIRE_87 | SYNTHESIZED_WIRE_88;

assign	SYNTHESIZED_WIRE_58 = SYNTHESIZED_WIRE_81 | SYNTHESIZED_WIRE_89 | SYNTHESIZED_WIRE_90 | SYNTHESIZED_WIRE_82;

assign	SYNTHESIZED_WIRE_15 = SYNTHESIZED_WIRE_89 | SYNTHESIZED_WIRE_90 | SYNTHESIZED_WIRE_88;

assign	SYNTHESIZED_WIRE_16 = SYNTHESIZED_WIRE_89 | SYNTHESIZED_WIRE_87 | SYNTHESIZED_WIRE_91;

assign	SYNTHESIZED_WIRE_17 = SYNTHESIZED_WIRE_88 | SYNTHESIZED_WIRE_90 | SYNTHESIZED_WIRE_91;

assign	Sb = SYNTHESIZED_WIRE_15 & SYNTHESIZED_WIRE_16 & SYNTHESIZED_WIRE_17 & SYNTHESIZED_WIRE_18;

assign	SYNTHESIZED_WIRE_59 = SYNTHESIZED_WIRE_88 | SYNTHESIZED_WIRE_90 | SYNTHESIZED_WIRE_91;

assign	SYNTHESIZED_WIRE_60 = SYNTHESIZED_WIRE_88 | SYNTHESIZED_WIRE_89 | SYNTHESIZED_WIRE_91;

assign	SYNTHESIZED_WIRE_89 =  ~SYNTHESIZED_WIRE_86;

assign	SYNTHESIZED_WIRE_61 = SYNTHESIZED_WIRE_89 | SYNTHESIZED_WIRE_87 | SYNTHESIZED_WIRE_88;

assign	SYNTHESIZED_WIRE_62 = SYNTHESIZED_WIRE_81 | SYNTHESIZED_WIRE_86 | SYNTHESIZED_WIRE_87 | SYNTHESIZED_WIRE_82;

assign	SYNTHESIZED_WIRE_63 = SYNTHESIZED_WIRE_81 | SYNTHESIZED_WIRE_86 | SYNTHESIZED_WIRE_90 | SYNTHESIZED_WIRE_88;

assign	SYNTHESIZED_WIRE_64 = SYNTHESIZED_WIRE_91 | SYNTHESIZED_WIRE_89 | SYNTHESIZED_WIRE_90 | SYNTHESIZED_WIRE_82;

assign	SYNTHESIZED_WIRE_56 = SYNTHESIZED_WIRE_86 | SYNTHESIZED_WIRE_87 | SYNTHESIZED_WIRE_82;

assign	SYNTHESIZED_WIRE_57 = SYNTHESIZED_WIRE_88 | SYNTHESIZED_WIRE_86 | SYNTHESIZED_WIRE_81;

assign	SYNTHESIZED_WIRE_55 = SYNTHESIZED_WIRE_87 | SYNTHESIZED_WIRE_81;

assign	SYNTHESIZED_WIRE_65 = SYNTHESIZED_WIRE_82 | SYNTHESIZED_WIRE_87 | SYNTHESIZED_WIRE_81;

assign	SYNTHESIZED_WIRE_66 = SYNTHESIZED_WIRE_82 | SYNTHESIZED_WIRE_89 | SYNTHESIZED_WIRE_81;

assign	SYNTHESIZED_WIRE_67 = SYNTHESIZED_WIRE_89 | SYNTHESIZED_WIRE_87 | SYNTHESIZED_WIRE_81;

assign	SYNTHESIZED_WIRE_87 =  ~SYNTHESIZED_WIRE_90;

assign	SYNTHESIZED_WIRE_68 = SYNTHESIZED_WIRE_91 | SYNTHESIZED_WIRE_86 | SYNTHESIZED_WIRE_87 | SYNTHESIZED_WIRE_88;

assign	SYNTHESIZED_WIRE_53 = SYNTHESIZED_WIRE_81 | SYNTHESIZED_WIRE_89 | SYNTHESIZED_WIRE_87 | SYNTHESIZED_WIRE_88;

assign	SYNTHESIZED_WIRE_54 = SYNTHESIZED_WIRE_91 | SYNTHESIZED_WIRE_86 | SYNTHESIZED_WIRE_90 | SYNTHESIZED_WIRE_88;


always@(posedge SYNTHESIZED_WIRE_85 or negedge Reset or negedge SYNTHESIZED_WIRE_84)
begin
if (!Reset)
	begin
	SYNTHESIZED_WIRE_86 <= 0;
	end
else
if (!SYNTHESIZED_WIRE_84)
	begin
	SYNTHESIZED_WIRE_86 <= 1;
	end
else
	begin
	SYNTHESIZED_WIRE_86 <= SYNTHESIZED_WIRE_92;
	end
end

assign	SYNTHESIZED_WIRE_52 = SYNTHESIZED_WIRE_82 | SYNTHESIZED_WIRE_86 | SYNTHESIZED_WIRE_81;


always@(posedge SYNTHESIZED_WIRE_92 or negedge Reset or negedge SYNTHESIZED_WIRE_84)
begin
if (!Reset)
	begin
	SYNTHESIZED_WIRE_82 <= 0;
	end
else
if (!SYNTHESIZED_WIRE_84)
	begin
	SYNTHESIZED_WIRE_82 <= 1;
	end
else
	begin
	SYNTHESIZED_WIRE_82 <= SYNTHESIZED_WIRE_83;
	end
end

assign	SYNTHESIZED_WIRE_1 =  ~SYNTHESIZED_WIRE_81;

assign	SYNTHESIZED_WIRE_83 =  ~SYNTHESIZED_WIRE_82;

assign	SYNTHESIZED_WIRE_85 =  ~SYNTHESIZED_WIRE_90;

assign	Sg = SYNTHESIZED_WIRE_52 & SYNTHESIZED_WIRE_53 & SYNTHESIZED_WIRE_54;

assign	Se = SYNTHESIZED_WIRE_55 & SYNTHESIZED_WIRE_56 & SYNTHESIZED_WIRE_57;

assign	Sc = SYNTHESIZED_WIRE_58 & SYNTHESIZED_WIRE_59 & SYNTHESIZED_WIRE_60;

assign	Sd = SYNTHESIZED_WIRE_61 & SYNTHESIZED_WIRE_62 & SYNTHESIZED_WIRE_63 & SYNTHESIZED_WIRE_64;

assign	Sf = SYNTHESIZED_WIRE_65 & SYNTHESIZED_WIRE_66 & SYNTHESIZED_WIRE_67 & SYNTHESIZED_WIRE_68;

assign	SYNTHESIZED_WIRE_92 =  ~SYNTHESIZED_WIRE_86;


assign	SYNTHESIZED_WIRE_77 = SYNTHESIZED_WIRE_81 | SYNTHESIZED_WIRE_86 | SYNTHESIZED_WIRE_87 | SYNTHESIZED_WIRE_82;

assign	SYNTHESIZED_WIRE_78 = SYNTHESIZED_WIRE_81 | SYNTHESIZED_WIRE_86 | SYNTHESIZED_WIRE_90 | SYNTHESIZED_WIRE_88;

assign	SYNTHESIZED_WIRE_79 = SYNTHESIZED_WIRE_91 | SYNTHESIZED_WIRE_89 | SYNTHESIZED_WIRE_87 | SYNTHESIZED_WIRE_82;

assign	SYNTHESIZED_WIRE_80 = SYNTHESIZED_WIRE_91 | SYNTHESIZED_WIRE_86 | SYNTHESIZED_WIRE_87 | SYNTHESIZED_WIRE_88;

assign	Sa = SYNTHESIZED_WIRE_77 & SYNTHESIZED_WIRE_78 & SYNTHESIZED_WIRE_79 & SYNTHESIZED_WIRE_80;


endmodule
